`timescale 1ns / 1ps

module de_compress_flag(
	
    );
endmodule
